library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

entity ram_512x8 is
    Port ( 
		  clk		: in  std_logic;
        reset	: in  std_logic;
        Din		: in  std_logic_vector(7 downto 0);
        WrEn	: in  std_logic;
        RdEn	: in  std_logic;
        Dout	: out std_logic_vector(7 downto 0);
		  RdAddr : in  std_logic_vector(12 downto 0)
	);
end ram_512x8;

architecture Behavioral of ram_512x8 is	
	type ram_type is array (0 to 8191) of std_logic_vector (7 downto 0);
	signal RAM 			: ram_type := (  
												x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"4D",x"41",x"49",x"4E",x"20",x"4D",x"45",x"4E",x"55",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"0A",
												x"20",x"20",x"20",x"20",x"20",x"20",x"28",x"31",x"29",x"53",x"74",x"61",x"6E",x"64",x"61",x"72",x"64",x"20",x"4D",x"6F",x"64",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"0A",
												x"20",x"20",x"20",x"20",x"20",x"20",x"28",x"32",x"29",x"52",x"61",x"73",x"74",x"67",x"65",x"6C",x"65",x"20",x"4D",x"6F",x"64",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"0A",
												x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"28",x"33",x"29",x"50",x"52",x"42",x"53",x"20",x"4D",x"6F",x"64",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"0A",
												x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"0A",
												x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"0A",
												x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"0A",
												x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"0A",
												
												x"20",x"20",x"20",x"20",x"28",x"31",x"29",x"46",x"72",x"65",x"71",x"75",x"65",x"6E",x"63",x"79",x"20",x"56",x"61",x"6C",x"75",x"65",x"73",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"0A",
												x"20",x"20",x"20",x"20",x"20",x"28",x"32",x"29",x"53",x"74",x"65",x"70",x"53",x"69",x"7A",x"65",x"20",x"56",x"61",x"6C",x"75",x"65",x"73",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"0A",
												x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"0A",
												x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"0A",
												x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"0A",
												x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"0A",
												x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"0A",
												x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"0A",
												
												x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"46",x"72",x"65",x"71",x"75",x"65",x"6E",x"63",x"79",x"20",x"56",x"61",x"6C",x"75",x"65",x"73",x"20",x"20",x"20",x"20",x"20",x"20",x"0A",
												x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"33",x"32",x"20",x"64",x"69",x"67",x"69",x"74",x"20",x"62",x"65",x"67",x"69",x"6E",x"6E",x"69",x"6E",x"67",x"20",x"20",x"20",x"20",x"20",x"0A",
												x"20",x"20",x"20",x"66",x"72",x"6F",x"6D",x"20",x"74",x"68",x"65",x"20",x"6C",x"6F",x"77",x"65",x"73",x"74",x"20",x"66",x"72",x"65",x"71",x"75",x"65",x"6E",x"63",x"79",x"20",x"20",x"20",x"0A",
												x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"0A",
												x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"0A",
												x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"0A",
												x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"0A",
												x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"0A",
												
												x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"53",x"74",x"65",x"70",x"53",x"69",x"7A",x"65",x"20",x"56",x"61",x"6C",x"75",x"65",x"73",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"0A",
												x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"33",x"20",x"64",x"69",x"67",x"69",x"74",x"20",x"66",x"6F",x"72",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"0A",
												x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"31",x"20",x"53",x"74",x"65",x"70",x"20",x"53",x"69",x"7A",x"65",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"0A",
												x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"0A",
												x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"0A",
												x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"0A",
												x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"0A",
												x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"0A",
												
												x"20",x"20",x"20",x"20",x"28",x"31",x"29",x"46",x"72",x"65",x"71",x"75",x"65",x"6E",x"63",x"79",x"20",x"56",x"61",x"6C",x"75",x"65",x"73",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"0A",
												x"20",x"20",x"20",x"20",x"20",x"28",x"32",x"29",x"53",x"74",x"65",x"70",x"53",x"69",x"7A",x"65",x"20",x"56",x"61",x"6C",x"75",x"65",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"0A",
												x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"0A",
												x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"0A",
												x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"0A",
												x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"0A",
												x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"0A",
												x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"0A",
												
												x"20",x"20",x"20",x"20",x"46",x"72",x"65",x"71",x"75",x"65",x"6E",x"63",x"79",x"20",x"56",x"61",x"6C",x"75",x"65",x"73",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"0A",
												x"20",x"20",x"33",x"32",x"20",x"44",x"69",x"67",x"69",x"74",x"73",x"20",x"66",x"72",x"6F",x"6D",x"20",x"74",x"68",x"65",x"20",x"6C",x"6F",x"77",x"65",x"73",x"74",x"20",x"20",x"20",x"20",x"0A",
												x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"0A",
												x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"0A",
												x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"0A",
												x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"0A",
												x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"0A",
												x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"0A",
												
												x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"53",x"74",x"65",x"70",x"53",x"69",x"7A",x"65",x"20",x"56",x"61",x"6C",x"75",x"65",x"73",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"0A",
												x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"33",x"20",x"64",x"69",x"67",x"69",x"74",x"20",x"66",x"6F",x"72",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"0A",
												x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"31",x"20",x"53",x"74",x"65",x"70",x"20",x"53",x"69",x"7A",x"65",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"0A",
												x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"0A",
												x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"0A",
												x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"0A",
												x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"0A",
												x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"0A",
												
												x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"28",x"31",x"29",x"4D",x"65",x"72",x"6B",x"65",x"7A",x"20",x"46",x"72",x"65",x"6B",x"61",x"6E",x"73",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"0A",
												x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"28",x"32",x"29",x"46",x"72",x"65",x"6B",x"61",x"6E",x"73",x"20",x"42",x"61",x"6E",x"64",x"69",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"0A",
												x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"0A",
												x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"0A",
												x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"0A",
												x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"0A",
												x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"0A",
												x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"0A",
												
												x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"4D",x"65",x"72",x"6B",x"65",x"7A",x"20",x"46",x"72",x"65",x"6B",x"61",x"6E",x"73",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"0A",
												x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"38",x"20",x"44",x"69",x"67",x"69",x"74",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"0A",
												x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"0A",
												x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"0A",
												x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"0A",
												x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"0A",
												x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"0A",
												x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"0A",
												
												x"31",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"46",x"72",x"65",x"6B",x"61",x"6E",x"73",x"20",x"42",x"61",x"6E",x"64",x"69",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"0A",
												x"31",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"38",x"20",x"44",x"69",x"67",x"69",x"74",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"0A",
												x"31",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"0A",
												x"31",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"0A",
												x"31",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"0A",
												x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"0A",
												x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"0A",
												x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"0A",
		 
												
												x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"28",x"31",x"29",x"31",x"2E",x"42",x"61",x"6E",x"74",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"0A",
												x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"28",x"32",x"29",x"32",x"2E",x"42",x"61",x"6E",x"74",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"0A",
												x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"28",x"33",x"29",x"33",x"2E",x"42",x"61",x"6E",x"74",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"0A",
												x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"28",x"34",x"29",x"34",x"2E",x"42",x"61",x"6E",x"74",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"0A",
												x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"0A",
												x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"0A",
												x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"0A",
												x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"0A",
												
												x"52",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"50",x"4F",x"57",x"45",x"52",x"20",x"50",x"52",x"4F",x"46",x"49",x"4C",x"45",x"31",x"20",x"20",x"20",x"20",x"20",x"0A",
												x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"50",x"4F",x"57",x"45",x"52",x"20",x"50",x"52",x"4F",x"46",x"49",x"4C",x"45",x"32",x"20",x"20",x"20",x"20",x"20",x"0A",
												x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"50",x"4F",x"57",x"45",x"52",x"20",x"50",x"52",x"4F",x"46",x"49",x"4C",x"45",x"33",x"20",x"20",x"20",x"20",x"20",x"0A",
												x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"50",x"4F",x"57",x"45",x"52",x"20",x"50",x"52",x"4F",x"46",x"49",x"4C",x"45",x"34",x"20",x"20",x"20",x"20",x"20",x"0A",
												x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"50",x"4F",x"57",x"45",x"52",x"20",x"50",x"52",x"4F",x"46",x"49",x"4C",x"45",x"35",x"20",x"20",x"20",x"20",x"20",x"0A",
												x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"50",x"4F",x"57",x"45",x"52",x"20",x"50",x"52",x"4F",x"46",x"49",x"4C",x"45",x"36",x"20",x"20",x"20",x"20",x"20",x"0A",
												x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"50",x"4F",x"57",x"45",x"52",x"20",x"50",x"52",x"4F",x"46",x"49",x"4C",x"45",x"37",x"20",x"20",x"20",x"20",x"20",x"0A",
												x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"50",x"4F",x"57",x"45",x"52",x"20",x"50",x"52",x"4F",x"46",x"49",x"4C",x"45",x"38",x"20",x"20",x"20",x"20",x"20",x"0A",
												
												x"49",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"4F",x"50",x"54",x"49",x"53",x"49",x"53",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"0A",
												x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"4E",x"45",x"57",x"20",x"4D",x"45",x"4E",x"55",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"0A",
												x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"41",x"4C",x"54",x"20",x"4D",x"45",x"4E",x"55",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"0A",
												x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"4F",x"50",x"54",x"49",x"4F",x"4E",x"53",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"0A",
												x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"43",x"52",x"45",x"44",x"49",x"54",x"53",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"0A",
												x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"50",x"52",x"4F",x"4A",x"45",x"43",x"54",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"0A",
												x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"52",x"41",x"4D",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"0A",
												x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"54",x"52",x"41",x"4E",x"53",x"4D",x"49",x"54",x"54",x"45",x"52",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"0A",
												
												x"50",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"42",x"41",x"55",x"44",x"20",x"46",x"52",x"45",x"51",x"55",x"45",x"4E",x"43",x"49",x"45",x"53",x"20",x"20",x"20",x"20",x"20",x"0A",
												x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"42",x"41",x"55",x"44",x"32",x"20",x"46",x"52",x"45",x"51",x"55",x"45",x"4E",x"43",x"49",x"45",x"53",x"20",x"20",x"20",x"20",x"0A",
												x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"42",x"41",x"55",x"44",x"33",x"20",x"46",x"52",x"45",x"51",x"55",x"45",x"4E",x"43",x"49",x"45",x"53",x"20",x"20",x"20",x"20",x"0A",
												x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"42",x"41",x"55",x"44",x"34",x"20",x"46",x"52",x"45",x"51",x"55",x"45",x"4E",x"43",x"49",x"45",x"53",x"20",x"20",x"20",x"20",x"0A",
												x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"42",x"41",x"55",x"44",x"35",x"20",x"46",x"52",x"45",x"51",x"55",x"45",x"4E",x"43",x"49",x"45",x"53",x"20",x"20",x"20",x"20",x"0A",
												x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"42",x"41",x"55",x"44",x"36",x"20",x"46",x"52",x"45",x"51",x"55",x"45",x"4E",x"43",x"49",x"45",x"53",x"20",x"20",x"20",x"20",x"0A",
												x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"42",x"41",x"55",x"44",x"37",x"20",x"46",x"52",x"45",x"51",x"55",x"45",x"4E",x"43",x"49",x"45",x"53",x"20",x"20",x"20",x"20",x"0A",
												x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"42",x"41",x"55",x"44",x"38",x"20",x"46",x"52",x"45",x"51",x"55",x"45",x"4E",x"43",x"49",x"45",x"53",x"20",x"20",x"20",x"20",x"0A",
												
												x"51",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"53",x"57",x"45",x"45",x"50",x"20",x"56",x"45",x"4C",x"4F",x"43",x"49",x"54",x"59",x"31",x"20",x"20",x"20",x"20",x"0A",
												x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"53",x"57",x"45",x"45",x"50",x"20",x"56",x"45",x"4C",x"4F",x"43",x"49",x"54",x"59",x"32",x"20",x"20",x"20",x"20",x"0A",
												x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"53",x"57",x"45",x"45",x"50",x"20",x"56",x"45",x"4C",x"4F",x"43",x"49",x"54",x"59",x"33",x"20",x"20",x"20",x"20",x"0A",
												x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"53",x"57",x"45",x"45",x"50",x"20",x"56",x"45",x"4C",x"4F",x"43",x"49",x"54",x"59",x"34",x"20",x"20",x"20",x"20",x"0A",
												x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"53",x"57",x"45",x"45",x"50",x"20",x"56",x"45",x"4C",x"4F",x"43",x"49",x"54",x"59",x"35",x"20",x"20",x"20",x"20",x"0A",
												x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"53",x"57",x"45",x"45",x"50",x"20",x"56",x"45",x"4C",x"4F",x"43",x"49",x"54",x"59",x"36",x"20",x"20",x"20",x"20",x"0A",
												x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"53",x"57",x"45",x"45",x"50",x"20",x"56",x"45",x"4C",x"4F",x"43",x"49",x"54",x"59",x"37",x"20",x"20",x"20",x"20",x"0A",
												x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"53",x"57",x"45",x"45",x"50",x"20",x"56",x"45",x"4C",x"4F",x"43",x"49",x"54",x"59",x"38",x"20",x"20",x"20",x"20",x"0A",
												
												x"52",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"50",x"4F",x"57",x"45",x"52",x"20",x"50",x"52",x"4F",x"46",x"49",x"4C",x"45",x"31",x"20",x"20",x"20",x"20",x"20",x"0A",
												x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"50",x"4F",x"57",x"45",x"52",x"20",x"50",x"52",x"4F",x"46",x"49",x"4C",x"45",x"32",x"20",x"20",x"20",x"20",x"20",x"0A",
												x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"50",x"4F",x"57",x"45",x"52",x"20",x"50",x"52",x"4F",x"46",x"49",x"4C",x"45",x"33",x"20",x"20",x"20",x"20",x"20",x"0A",
												x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"50",x"4F",x"57",x"45",x"52",x"20",x"50",x"52",x"4F",x"46",x"49",x"4C",x"45",x"34",x"20",x"20",x"20",x"20",x"20",x"0A",
												x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"50",x"4F",x"57",x"45",x"52",x"20",x"50",x"52",x"4F",x"46",x"49",x"4C",x"45",x"35",x"20",x"20",x"20",x"20",x"20",x"0A",
												x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"50",x"4F",x"57",x"45",x"52",x"20",x"50",x"52",x"4F",x"46",x"49",x"4C",x"45",x"36",x"20",x"20",x"20",x"20",x"20",x"0A",
												x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"50",x"4F",x"57",x"45",x"52",x"20",x"50",x"52",x"4F",x"46",x"49",x"4C",x"45",x"37",x"20",x"20",x"20",x"20",x"20",x"0A",
												x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"50",x"4F",x"57",x"45",x"52",x"20",x"50",x"52",x"4F",x"46",x"49",x"4C",x"45",x"38",x"20",x"20",x"20",x"20",x"20",x"0A",
												
												x"49",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"4F",x"50",x"54",x"49",x"53",x"49",x"53",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"0A",
												x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"4E",x"45",x"57",x"20",x"4D",x"45",x"4E",x"55",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"0A",
												x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"41",x"4C",x"54",x"20",x"4D",x"45",x"4E",x"55",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"0A",
												x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"4F",x"50",x"54",x"49",x"4F",x"4E",x"53",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"0A",
												x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"43",x"52",x"45",x"44",x"49",x"54",x"53",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"0A",
												x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"50",x"52",x"4F",x"4A",x"45",x"43",x"54",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"0A",
												x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"52",x"41",x"4D",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"0A",
												x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"54",x"52",x"41",x"4E",x"53",x"4D",x"49",x"54",x"54",x"45",x"52",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"0A",
												
												x"50",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"42",x"41",x"55",x"44",x"20",x"46",x"52",x"45",x"51",x"55",x"45",x"4E",x"43",x"49",x"45",x"53",x"20",x"20",x"20",x"20",x"20",x"0A",
												x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"42",x"41",x"55",x"44",x"32",x"20",x"46",x"52",x"45",x"51",x"55",x"45",x"4E",x"43",x"49",x"45",x"53",x"20",x"20",x"20",x"20",x"0A",
												x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"42",x"41",x"55",x"44",x"33",x"20",x"46",x"52",x"45",x"51",x"55",x"45",x"4E",x"43",x"49",x"45",x"53",x"20",x"20",x"20",x"20",x"0A",
												x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"42",x"41",x"55",x"44",x"34",x"20",x"46",x"52",x"45",x"51",x"55",x"45",x"4E",x"43",x"49",x"45",x"53",x"20",x"20",x"20",x"20",x"0A",
												x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"42",x"41",x"55",x"44",x"35",x"20",x"46",x"52",x"45",x"51",x"55",x"45",x"4E",x"43",x"49",x"45",x"53",x"20",x"20",x"20",x"20",x"0A",
												x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"42",x"41",x"55",x"44",x"36",x"20",x"46",x"52",x"45",x"51",x"55",x"45",x"4E",x"43",x"49",x"45",x"53",x"20",x"20",x"20",x"20",x"0A",
												x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"42",x"41",x"55",x"44",x"37",x"20",x"46",x"52",x"45",x"51",x"55",x"45",x"4E",x"43",x"49",x"45",x"53",x"20",x"20",x"20",x"20",x"0A",
												x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"42",x"41",x"55",x"44",x"38",x"20",x"46",x"52",x"45",x"51",x"55",x"45",x"4E",x"43",x"49",x"45",x"53",x"20",x"20",x"20",x"20",x"0A",
												
												x"51",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"53",x"57",x"45",x"45",x"50",x"20",x"56",x"45",x"4C",x"4F",x"43",x"49",x"54",x"59",x"31",x"20",x"20",x"20",x"20",x"0A",
												x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"53",x"57",x"45",x"45",x"50",x"20",x"56",x"45",x"4C",x"4F",x"43",x"49",x"54",x"59",x"32",x"20",x"20",x"20",x"20",x"0A",
												x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"53",x"57",x"45",x"45",x"50",x"20",x"56",x"45",x"4C",x"4F",x"43",x"49",x"54",x"59",x"33",x"20",x"20",x"20",x"20",x"0A",
												x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"53",x"57",x"45",x"45",x"50",x"20",x"56",x"45",x"4C",x"4F",x"43",x"49",x"54",x"59",x"34",x"20",x"20",x"20",x"20",x"0A",
												x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"53",x"57",x"45",x"45",x"50",x"20",x"56",x"45",x"4C",x"4F",x"43",x"49",x"54",x"59",x"35",x"20",x"20",x"20",x"20",x"0A",
												x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"53",x"57",x"45",x"45",x"50",x"20",x"56",x"45",x"4C",x"4F",x"43",x"49",x"54",x"59",x"36",x"20",x"20",x"20",x"20",x"0A",
												x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"53",x"57",x"45",x"45",x"50",x"20",x"56",x"45",x"4C",x"4F",x"43",x"49",x"54",x"59",x"37",x"20",x"20",x"20",x"20",x"0A",
												x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"53",x"57",x"45",x"45",x"50",x"20",x"56",x"45",x"4C",x"4F",x"43",x"49",x"54",x"59",x"38",x"20",x"20",x"20",x"20",x"0A",
												
												x"52",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"50",x"4F",x"57",x"45",x"52",x"20",x"50",x"52",x"4F",x"46",x"49",x"4C",x"45",x"31",x"20",x"20",x"20",x"20",x"20",x"0A",
												x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"50",x"4F",x"57",x"45",x"52",x"20",x"50",x"52",x"4F",x"46",x"49",x"4C",x"45",x"32",x"20",x"20",x"20",x"20",x"20",x"0A",
												x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"50",x"4F",x"57",x"45",x"52",x"20",x"50",x"52",x"4F",x"46",x"49",x"4C",x"45",x"33",x"20",x"20",x"20",x"20",x"20",x"0A",
												x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"50",x"4F",x"57",x"45",x"52",x"20",x"50",x"52",x"4F",x"46",x"49",x"4C",x"45",x"34",x"20",x"20",x"20",x"20",x"20",x"0A",
												x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"50",x"4F",x"57",x"45",x"52",x"20",x"50",x"52",x"4F",x"46",x"49",x"4C",x"45",x"35",x"20",x"20",x"20",x"20",x"20",x"0A",
												x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"50",x"4F",x"57",x"45",x"52",x"20",x"50",x"52",x"4F",x"46",x"49",x"4C",x"45",x"36",x"20",x"20",x"20",x"20",x"20",x"0A",
												x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"50",x"4F",x"57",x"45",x"52",x"20",x"50",x"52",x"4F",x"46",x"49",x"4C",x"45",x"37",x"20",x"20",x"20",x"20",x"20",x"0A",
												x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"50",x"4F",x"57",x"45",x"52",x"20",x"50",x"52",x"4F",x"46",x"49",x"4C",x"45",x"38",x"20",x"20",x"20",x"20",x"20",x"0A",
												
												x"49",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"4F",x"50",x"54",x"49",x"53",x"49",x"53",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"0A",
												x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"4E",x"45",x"57",x"20",x"4D",x"45",x"4E",x"55",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"0A",
												x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"41",x"4C",x"54",x"20",x"4D",x"45",x"4E",x"55",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"0A",
												x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"4F",x"50",x"54",x"49",x"4F",x"4E",x"53",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"0A",
												x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"43",x"52",x"45",x"44",x"49",x"54",x"53",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"0A",
												x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"50",x"52",x"4F",x"4A",x"45",x"43",x"54",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"0A",
												x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"52",x"41",x"4D",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"0A",
												x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"54",x"52",x"41",x"4E",x"53",x"4D",x"49",x"54",x"54",x"45",x"52",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"0A",
												
												x"50",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"42",x"41",x"55",x"44",x"20",x"46",x"52",x"45",x"51",x"55",x"45",x"4E",x"43",x"49",x"45",x"53",x"20",x"20",x"20",x"20",x"20",x"0A",
												x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"42",x"41",x"55",x"44",x"32",x"20",x"46",x"52",x"45",x"51",x"55",x"45",x"4E",x"43",x"49",x"45",x"53",x"20",x"20",x"20",x"20",x"0A",
												x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"42",x"41",x"55",x"44",x"33",x"20",x"46",x"52",x"45",x"51",x"55",x"45",x"4E",x"43",x"49",x"45",x"53",x"20",x"20",x"20",x"20",x"0A",
												x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"42",x"41",x"55",x"44",x"34",x"20",x"46",x"52",x"45",x"51",x"55",x"45",x"4E",x"43",x"49",x"45",x"53",x"20",x"20",x"20",x"20",x"0A",
												x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"42",x"41",x"55",x"44",x"35",x"20",x"46",x"52",x"45",x"51",x"55",x"45",x"4E",x"43",x"49",x"45",x"53",x"20",x"20",x"20",x"20",x"0A",
												x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"42",x"41",x"55",x"44",x"36",x"20",x"46",x"52",x"45",x"51",x"55",x"45",x"4E",x"43",x"49",x"45",x"53",x"20",x"20",x"20",x"20",x"0A",
												x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"42",x"41",x"55",x"44",x"37",x"20",x"46",x"52",x"45",x"51",x"55",x"45",x"4E",x"43",x"49",x"45",x"53",x"20",x"20",x"20",x"20",x"0A",
												x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"42",x"41",x"55",x"44",x"38",x"20",x"46",x"52",x"45",x"51",x"55",x"45",x"4E",x"43",x"49",x"45",x"53",x"20",x"20",x"20",x"20",x"0A",
												
												x"51",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"53",x"57",x"45",x"45",x"50",x"20",x"56",x"45",x"4C",x"4F",x"43",x"49",x"54",x"59",x"31",x"20",x"20",x"20",x"20",x"0A",
												x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"53",x"57",x"45",x"45",x"50",x"20",x"56",x"45",x"4C",x"4F",x"43",x"49",x"54",x"59",x"32",x"20",x"20",x"20",x"20",x"0A",
												x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"53",x"57",x"45",x"45",x"50",x"20",x"56",x"45",x"4C",x"4F",x"43",x"49",x"54",x"59",x"33",x"20",x"20",x"20",x"20",x"0A",
												x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"53",x"57",x"45",x"45",x"50",x"20",x"56",x"45",x"4C",x"4F",x"43",x"49",x"54",x"59",x"34",x"20",x"20",x"20",x"20",x"0A",
												x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"53",x"57",x"45",x"45",x"50",x"20",x"56",x"45",x"4C",x"4F",x"43",x"49",x"54",x"59",x"35",x"20",x"20",x"20",x"20",x"0A",
												x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"53",x"57",x"45",x"45",x"50",x"20",x"56",x"45",x"4C",x"4F",x"43",x"49",x"54",x"59",x"36",x"20",x"20",x"20",x"20",x"0A",
												x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"53",x"57",x"45",x"45",x"50",x"20",x"56",x"45",x"4C",x"4F",x"43",x"49",x"54",x"59",x"37",x"20",x"20",x"20",x"20",x"0A",
												x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"53",x"57",x"45",x"45",x"50",x"20",x"56",x"45",x"4C",x"4F",x"43",x"49",x"54",x"59",x"38",x"20",x"20",x"20",x"20",x"0A",
												
												x"52",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"50",x"4F",x"57",x"45",x"52",x"20",x"50",x"52",x"4F",x"46",x"49",x"4C",x"45",x"31",x"20",x"20",x"20",x"20",x"20",x"0A",
												x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"50",x"4F",x"57",x"45",x"52",x"20",x"50",x"52",x"4F",x"46",x"49",x"4C",x"45",x"32",x"20",x"20",x"20",x"20",x"20",x"0A",
												x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"50",x"4F",x"57",x"45",x"52",x"20",x"50",x"52",x"4F",x"46",x"49",x"4C",x"45",x"33",x"20",x"20",x"20",x"20",x"20",x"0A",
												x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"50",x"4F",x"57",x"45",x"52",x"20",x"50",x"52",x"4F",x"46",x"49",x"4C",x"45",x"34",x"20",x"20",x"20",x"20",x"20",x"0A",
												x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"50",x"4F",x"57",x"45",x"52",x"20",x"50",x"52",x"4F",x"46",x"49",x"4C",x"45",x"35",x"20",x"20",x"20",x"20",x"20",x"0A",
												x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"50",x"4F",x"57",x"45",x"52",x"20",x"50",x"52",x"4F",x"46",x"49",x"4C",x"45",x"36",x"20",x"20",x"20",x"20",x"20",x"0A",
												x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"50",x"4F",x"57",x"45",x"52",x"20",x"50",x"52",x"4F",x"46",x"49",x"4C",x"45",x"37",x"20",x"20",x"20",x"20",x"20",x"0A",
												x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"50",x"4F",x"57",x"45",x"52",x"20",x"50",x"52",x"4F",x"46",x"49",x"4C",x"45",x"38",x"20",x"20",x"20",x"20",x"20",x"0A",
												
												x"49",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"4F",x"50",x"54",x"49",x"53",x"49",x"53",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"0A",
												x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"4E",x"45",x"57",x"20",x"4D",x"45",x"4E",x"55",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"0A",
												x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"41",x"4C",x"54",x"20",x"4D",x"45",x"4E",x"55",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"0A",
												x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"4F",x"50",x"54",x"49",x"4F",x"4E",x"53",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"0A",
												x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"43",x"52",x"45",x"44",x"49",x"54",x"53",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"0A",
												x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"50",x"52",x"4F",x"4A",x"45",x"43",x"54",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"0A",
												x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"52",x"41",x"4D",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"0A",
												x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"54",x"52",x"41",x"4E",x"53",x"4D",x"49",x"54",x"54",x"45",x"52",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"0A",
												
												x"50",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"42",x"41",x"55",x"44",x"20",x"46",x"52",x"45",x"51",x"55",x"45",x"4E",x"43",x"49",x"45",x"53",x"20",x"20",x"20",x"20",x"20",x"0A",
												x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"42",x"41",x"55",x"44",x"32",x"20",x"46",x"52",x"45",x"51",x"55",x"45",x"4E",x"43",x"49",x"45",x"53",x"20",x"20",x"20",x"20",x"0A",
												x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"42",x"41",x"55",x"44",x"33",x"20",x"46",x"52",x"45",x"51",x"55",x"45",x"4E",x"43",x"49",x"45",x"53",x"20",x"20",x"20",x"20",x"0A",
												x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"42",x"41",x"55",x"44",x"34",x"20",x"46",x"52",x"45",x"51",x"55",x"45",x"4E",x"43",x"49",x"45",x"53",x"20",x"20",x"20",x"20",x"0A",
												x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"42",x"41",x"55",x"44",x"35",x"20",x"46",x"52",x"45",x"51",x"55",x"45",x"4E",x"43",x"49",x"45",x"53",x"20",x"20",x"20",x"20",x"0A",
												x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"42",x"41",x"55",x"44",x"36",x"20",x"46",x"52",x"45",x"51",x"55",x"45",x"4E",x"43",x"49",x"45",x"53",x"20",x"20",x"20",x"20",x"0A",
												x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"42",x"41",x"55",x"44",x"37",x"20",x"46",x"52",x"45",x"51",x"55",x"45",x"4E",x"43",x"49",x"45",x"53",x"20",x"20",x"20",x"20",x"0A",
												x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"42",x"41",x"55",x"44",x"38",x"20",x"46",x"52",x"45",x"51",x"55",x"45",x"4E",x"43",x"49",x"45",x"53",x"20",x"20",x"20",x"20",x"0A",
												
												x"51",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"53",x"57",x"45",x"45",x"50",x"20",x"56",x"45",x"4C",x"4F",x"43",x"49",x"54",x"59",x"31",x"20",x"20",x"20",x"20",x"0A",
												x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"53",x"57",x"45",x"45",x"50",x"20",x"56",x"45",x"4C",x"4F",x"43",x"49",x"54",x"59",x"32",x"20",x"20",x"20",x"20",x"0A",
												x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"53",x"57",x"45",x"45",x"50",x"20",x"56",x"45",x"4C",x"4F",x"43",x"49",x"54",x"59",x"33",x"20",x"20",x"20",x"20",x"0A",
												x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"53",x"57",x"45",x"45",x"50",x"20",x"56",x"45",x"4C",x"4F",x"43",x"49",x"54",x"59",x"34",x"20",x"20",x"20",x"20",x"0A",
												x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"53",x"57",x"45",x"45",x"50",x"20",x"56",x"45",x"4C",x"4F",x"43",x"49",x"54",x"59",x"35",x"20",x"20",x"20",x"20",x"0A",
												x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"53",x"57",x"45",x"45",x"50",x"20",x"56",x"45",x"4C",x"4F",x"43",x"49",x"54",x"59",x"36",x"20",x"20",x"20",x"20",x"0A",
												x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"53",x"57",x"45",x"45",x"50",x"20",x"56",x"45",x"4C",x"4F",x"43",x"49",x"54",x"59",x"37",x"20",x"20",x"20",x"20",x"0A",
												x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"53",x"57",x"45",x"45",x"50",x"20",x"56",x"45",x"4C",x"4F",x"43",x"49",x"54",x"59",x"38",x"20",x"20",x"20",x"20",x"0A",
												
												x"52",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"50",x"4F",x"57",x"45",x"52",x"20",x"50",x"52",x"4F",x"46",x"49",x"4C",x"45",x"31",x"20",x"20",x"20",x"20",x"20",x"0A",
												x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"50",x"4F",x"57",x"45",x"52",x"20",x"50",x"52",x"4F",x"46",x"49",x"4C",x"45",x"32",x"20",x"20",x"20",x"20",x"20",x"0A",
												x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"50",x"4F",x"57",x"45",x"52",x"20",x"50",x"52",x"4F",x"46",x"49",x"4C",x"45",x"33",x"20",x"20",x"20",x"20",x"20",x"0A",
												x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"50",x"4F",x"57",x"45",x"52",x"20",x"50",x"52",x"4F",x"46",x"49",x"4C",x"45",x"34",x"20",x"20",x"20",x"20",x"20",x"0A",
												x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"50",x"4F",x"57",x"45",x"52",x"20",x"50",x"52",x"4F",x"46",x"49",x"4C",x"45",x"35",x"20",x"20",x"20",x"20",x"20",x"0A",
												x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"50",x"4F",x"57",x"45",x"52",x"20",x"50",x"52",x"4F",x"46",x"49",x"4C",x"45",x"36",x"20",x"20",x"20",x"20",x"20",x"0A",
												x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"50",x"4F",x"57",x"45",x"52",x"20",x"50",x"52",x"4F",x"46",x"49",x"4C",x"45",x"37",x"20",x"20",x"20",x"20",x"20",x"0A",
												x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"50",x"4F",x"57",x"45",x"52",x"20",x"50",x"52",x"4F",x"46",x"49",x"4C",x"45",x"38",x"20",x"20",x"20",x"20",x"20",x"0A",
												
												x"49",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"4F",x"50",x"54",x"49",x"53",x"49",x"53",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"0A",
												x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"4E",x"45",x"57",x"20",x"4D",x"45",x"4E",x"55",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"0A",
												x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"41",x"4C",x"54",x"20",x"4D",x"45",x"4E",x"55",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"0A",
												x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"4F",x"50",x"54",x"49",x"4F",x"4E",x"53",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"0A",
												x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"43",x"52",x"45",x"44",x"49",x"54",x"53",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"0A",
												x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"50",x"52",x"4F",x"4A",x"45",x"43",x"54",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"0A",
												x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"52",x"41",x"4D",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"0A",
												x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"54",x"52",x"41",x"4E",x"53",x"4D",x"49",x"54",x"54",x"45",x"52",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"0A",
												
												x"50",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"42",x"41",x"55",x"44",x"20",x"46",x"52",x"45",x"51",x"55",x"45",x"4E",x"43",x"49",x"45",x"53",x"20",x"20",x"20",x"20",x"20",x"0A",
												x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"42",x"41",x"55",x"44",x"32",x"20",x"46",x"52",x"45",x"51",x"55",x"45",x"4E",x"43",x"49",x"45",x"53",x"20",x"20",x"20",x"20",x"0A",
												x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"42",x"41",x"55",x"44",x"33",x"20",x"46",x"52",x"45",x"51",x"55",x"45",x"4E",x"43",x"49",x"45",x"53",x"20",x"20",x"20",x"20",x"0A",
												x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"42",x"41",x"55",x"44",x"34",x"20",x"46",x"52",x"45",x"51",x"55",x"45",x"4E",x"43",x"49",x"45",x"53",x"20",x"20",x"20",x"20",x"0A",
												x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"42",x"41",x"55",x"44",x"35",x"20",x"46",x"52",x"45",x"51",x"55",x"45",x"4E",x"43",x"49",x"45",x"53",x"20",x"20",x"20",x"20",x"0A",
												x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"42",x"41",x"55",x"44",x"36",x"20",x"46",x"52",x"45",x"51",x"55",x"45",x"4E",x"43",x"49",x"45",x"53",x"20",x"20",x"20",x"20",x"0A",
												x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"42",x"41",x"55",x"44",x"37",x"20",x"46",x"52",x"45",x"51",x"55",x"45",x"4E",x"43",x"49",x"45",x"53",x"20",x"20",x"20",x"20",x"0A",
												x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"42",x"41",x"55",x"44",x"38",x"20",x"46",x"52",x"45",x"51",x"55",x"45",x"4E",x"43",x"49",x"45",x"53",x"20",x"20",x"20",x"20",x"0A",
												
												x"51",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"53",x"57",x"45",x"45",x"50",x"20",x"56",x"45",x"4C",x"4F",x"43",x"49",x"54",x"59",x"31",x"20",x"20",x"20",x"20",x"0A",
												x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"53",x"57",x"45",x"45",x"50",x"20",x"56",x"45",x"4C",x"4F",x"43",x"49",x"54",x"59",x"32",x"20",x"20",x"20",x"20",x"0A",
												x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"53",x"57",x"45",x"45",x"50",x"20",x"56",x"45",x"4C",x"4F",x"43",x"49",x"54",x"59",x"33",x"20",x"20",x"20",x"20",x"0A",
												x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"53",x"57",x"45",x"45",x"50",x"20",x"56",x"45",x"4C",x"4F",x"43",x"49",x"54",x"59",x"34",x"20",x"20",x"20",x"20",x"0A",
												x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"53",x"57",x"45",x"45",x"50",x"20",x"56",x"45",x"4C",x"4F",x"43",x"49",x"54",x"59",x"35",x"20",x"20",x"20",x"20",x"0A",
												x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"53",x"57",x"45",x"45",x"50",x"20",x"56",x"45",x"4C",x"4F",x"43",x"49",x"54",x"59",x"36",x"20",x"20",x"20",x"20",x"0A",
												x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"53",x"57",x"45",x"45",x"50",x"20",x"56",x"45",x"4C",x"4F",x"43",x"49",x"54",x"59",x"37",x"20",x"20",x"20",x"20",x"0A",
												x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"53",x"57",x"45",x"45",x"50",x"20",x"56",x"45",x"4C",x"4F",x"43",x"49",x"54",x"59",x"38",x"20",x"20",x"20",x"20",x"0A",
												
												x"52",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"50",x"4F",x"57",x"45",x"52",x"20",x"50",x"52",x"4F",x"46",x"49",x"4C",x"45",x"31",x"20",x"20",x"20",x"20",x"20",x"0A",
												x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"50",x"4F",x"57",x"45",x"52",x"20",x"50",x"52",x"4F",x"46",x"49",x"4C",x"45",x"32",x"20",x"20",x"20",x"20",x"20",x"0A",
												x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"50",x"4F",x"57",x"45",x"52",x"20",x"50",x"52",x"4F",x"46",x"49",x"4C",x"45",x"33",x"20",x"20",x"20",x"20",x"20",x"0A",
												x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"50",x"4F",x"57",x"45",x"52",x"20",x"50",x"52",x"4F",x"46",x"49",x"4C",x"45",x"34",x"20",x"20",x"20",x"20",x"20",x"0A",
												x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"50",x"4F",x"57",x"45",x"52",x"20",x"50",x"52",x"4F",x"46",x"49",x"4C",x"45",x"35",x"20",x"20",x"20",x"20",x"20",x"0A",
												x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"50",x"4F",x"57",x"45",x"52",x"20",x"50",x"52",x"4F",x"46",x"49",x"4C",x"45",x"36",x"20",x"20",x"20",x"20",x"20",x"0A",
												x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"50",x"4F",x"57",x"45",x"52",x"20",x"50",x"52",x"4F",x"46",x"49",x"4C",x"45",x"37",x"20",x"20",x"20",x"20",x"20",x"0A",
												x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"50",x"4F",x"57",x"45",x"52",x"20",x"50",x"52",x"4F",x"46",x"49",x"4C",x"45",x"38",x"20",x"20",x"20",x"20",x"20",x"0A"
								); 
							
	
	signal WrAddr			: std_logic_vector(12 downto 0) := (others => '0');
	signal read_Address	: std_logic_vector(7 downto 0);
	
begin
	process (Clk,reset)
	begin
		if reset = '1' then
			WrAddr <= (others => '0');
		elsif rising_edge(Clk) then
			if WrEn = '1' then
				RAM(conv_integer(WrAddr)) <= Din;
				WrAddr <= WrAddr + '1';
			end if;
			
			if RdEn = '1' then
				Dout <= RAM(conv_integer(RdAddr));
			end if;
		end if;
	end process;
end Behavioral;